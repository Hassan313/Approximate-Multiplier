`timescale 1ns/1ns

module MULT_PPG16 (A, B, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);

input [15:0]A;
input [15:0]B;
output [15:0]PP0;
output [15:0]PP1;
output [15:0]PP2;
output [15:0]PP3;
output [15:0]PP4;
output [15:0]PP5;
output [15:0]PP6;
output [15:0]PP7;
output [15:0]PP8;
output [15:0]PP9;
output [15:0]PP10;
output [15:0]PP11;
output [15:0]PP12;
output [15:0]PP13;
output [15:0]PP14;
output [15:0]PP15;

////////////////// PP 0////////////////////////////
  AND2 U0 (.A1(A[0]),.A2(B[0]),.Z(PP0[0]));
  AND2 U1 (.A1(A[1]),.A2(B[0]),.Z(PP0[1]));
  AND2 U2 (.A1(A[2]),.A2(B[0]),.Z(PP0[2]));
  AND2 U3 (.A1(A[3]),.A2(B[0]),.Z(PP0[3]));
  AND2 U4 (.A1(A[4]),.A2(B[0]),.Z(PP0[4]));
  AND2 U5 (.A1(A[5]),.A2(B[0]),.Z(PP0[5]));
  AND2 U6 (.A1(A[6]),.A2(B[0]),.Z(PP0[6]));
  AND2 u7 (.A1(A[7]),.A2(B[0]),.Z(PP0[7]));
  AND2 UU0 (.A1(A[8]),.A2(B[0]),.Z(PP0[8]));
  AND2 UU1 (.A1(A[9]),.A2(B[0]),.Z(PP0[9]));
  AND2 UU2 (.A1(A[10]),.A2(B[0]),.Z(PP0[10]));
  AND2 UU3 (.A1(A[11]),.A2(B[0]),.Z(PP0[11]));
  AND2 UU4 (.A1(A[12]),.A2(B[0]),.Z(PP0[12]));
  AND2 UU5 (.A1(A[13]),.A2(B[0]),.Z(PP0[13]));
  AND2 UU6 (.A1(A[14]),.A2(B[0]),.Z(PP0[14]));
  AND2 uU7 (.A1(A[15]),.A2(B[0]),.Z(PP0[15]));
////////////////// PP 1////////////////////////////
  AND2 U7 (.A1(A[0]),.A2(B[1]),.Z(PP1[0]));
  AND2 U8 (.A1(A[1]),.A2(B[1]),.Z(PP1[1]));
  AND2 U9 (.A1(A[2]),.A2(B[1]),.Z(PP1[2]));
  AND2 U10 (.A1(A[3]),.A2(B[1]),.Z(PP1[3]));
  AND2 U11 (.A1(A[4]),.A2(B[1]),.Z(PP1[4]));
  AND2 U12 (.A1(A[5]),.A2(B[1]),.Z(PP1[5]));
  AND2 U13 (.A1(A[6]),.A2(B[1]),.Z(PP1[6]));
  AND2 u14 (.A1(A[7]),.A2(B[1]),.Z(PP1[7]));
  AND2 UU7 (.A1(A[8]),.A2(B[1]),.Z(PP1[8]));
  AND2 UU8 (.A1(A[9]),.A2(B[1]),.Z(PP1[9]));
  AND2 UU9 (.A1(A[10]),.A2(B[1]),.Z(PP1[10]));
  AND2 UU10 (.A1(A[11]),.A2(B[1]),.Z(PP1[11]));
  AND2 UU11 (.A1(A[12]),.A2(B[1]),.Z(PP1[12]));
  AND2 UU12 (.A1(A[13]),.A2(B[1]),.Z(PP1[13]));
  AND2 UU13 (.A1(A[14]),.A2(B[1]),.Z(PP1[14]));
  AND2 uU14 (.A1(A[15]),.A2(B[1]),.Z(PP1[15]));
////////////////// PP 2////////////////////////////
  AND2 U14 (.A1(A[0]),.A2(B[2]),.Z(PP2[0]));
  AND2 U15 (.A1(A[1]),.A2(B[2]),.Z(PP2[1]));
  AND2 U16 (.A1(A[2]),.A2(B[2]),.Z(PP2[2]));
  AND2 U17 (.A1(A[3]),.A2(B[2]),.Z(PP2[3]));
  AND2 U18 (.A1(A[4]),.A2(B[2]),.Z(PP2[4]));
  AND2 U19 (.A1(A[5]),.A2(B[2]),.Z(PP2[5]));
  AND2 U20 (.A1(A[6]),.A2(B[2]),.Z(PP2[6]));
  AND2 u21 (.A1(A[7]),.A2(B[2]),.Z(PP2[7]));
  AND2 UU14 (.A1(A[8]),.A2(B[2]),.Z(PP2[8]));
  AND2 UU15 (.A1(A[9]),.A2(B[2]),.Z(PP2[9]));
  AND2 UU16 (.A1(A[10]),.A2(B[2]),.Z(PP2[10]));
  AND2 UU17 (.A1(A[11]),.A2(B[2]),.Z(PP2[11]));
  AND2 UU18 (.A1(A[12]),.A2(B[2]),.Z(PP2[12]));
  AND2 UU19 (.A1(A[13]),.A2(B[2]),.Z(PP2[13]));
  AND2 UU20 (.A1(A[14]),.A2(B[2]),.Z(PP2[14]));
  AND2 Uu21 (.A1(A[15]),.A2(B[2]),.Z(PP2[15]));
////////////////// PP 3////////////////////////////
  AND2 U21 (.A1(A[0]),.A2(B[3]),.Z(PP3[0]));
  AND2 U22 (.A1(A[1]),.A2(B[3]),.Z(PP3[1]));
  AND2 U23 (.A1(A[2]),.A2(B[3]),.Z(PP3[2]));
  AND2 U24 (.A1(A[3]),.A2(B[3]),.Z(PP3[3]));
  AND2 U25 (.A1(A[4]),.A2(B[3]),.Z(PP3[4]));
  AND2 U26 (.A1(A[5]),.A2(B[3]),.Z(PP3[5]));
  AND2 U27 (.A1(A[6]),.A2(B[3]),.Z(PP3[6]));
  AND2 uU28 (.A1(A[7]),.A2(B[3]),.Z(PP3[7]));
  AND2 UU21 (.A1(A[8]),.A2(B[3]),.Z(PP3[8]));
  AND2 UU22 (.A1(A[9]),.A2(B[3]),.Z(PP3[9]));
  AND2 UU23 (.A1(A[10]),.A2(B[3]),.Z(PP3[10]));
  AND2 UU24 (.A1(A[11]),.A2(B[3]),.Z(PP3[11]));
  AND2 UU25 (.A1(A[12]),.A2(B[3]),.Z(PP3[12]));
  AND2 UU26 (.A1(A[13]),.A2(B[3]),.Z(PP3[13]));
  AND2 UU27 (.A1(A[14]),.A2(B[3]),.Z(PP3[14]));
  AND2 UT28 (.A1(A[15]),.A2(B[3]),.Z(PP3[15]));
////////////////// PP 4////////////////////////////
  AND2 U28 (.A1(A[0]),.A2(B[4]),.Z(PP4[0]));
  AND2 U29 (.A1(A[1]),.A2(B[4]),.Z(PP4[1]));
  AND2 U30 (.A1(A[2]),.A2(B[4]),.Z(PP4[2]));
  AND2 U31 (.A1(A[3]),.A2(B[4]),.Z(PP4[3]));
  AND2 U32 (.A1(A[4]),.A2(B[4]),.Z(PP4[4]));
  AND2 U33 (.A1(A[5]),.A2(B[4]),.Z(PP4[5]));
  AND2 U34 (.A1(A[6]),.A2(B[4]),.Z(PP4[6]));
  AND2 u35 (.A1(A[7]),.A2(B[4]),.Z(PP4[7]));
  AND2 UU28 (.A1(A[8]),.A2(B[4]),.Z(PP4[8]));
  AND2 UU29 (.A1(A[9]),.A2(B[4]),.Z(PP4[9]));
  AND2 UU30 (.A1(A[10]),.A2(B[4]),.Z(PP4[10]));
  AND2 UU31 (.A1(A[11]),.A2(B[4]),.Z(PP4[11]));
  AND2 UU32 (.A1(A[12]),.A2(B[4]),.Z(PP4[12]));
  AND2 UU33 (.A1(A[13]),.A2(B[4]),.Z(PP4[13]));
  AND2 UU34 (.A1(A[14]),.A2(B[4]),.Z(PP4[14]));
  AND2 uU35 (.A1(A[15]),.A2(B[4]),.Z(PP4[15]));
////////////////// PP 5////////////////////////////
  AND2 U35 (.A1(A[0]),.A2(B[5]),.Z(PP5[0]));
  AND2 U36 (.A1(A[1]),.A2(B[5]),.Z(PP5[1]));
  AND2 U37 (.A1(A[2]),.A2(B[5]),.Z(PP5[2]));
  AND2 U38 (.A1(A[3]),.A2(B[5]),.Z(PP5[3]));
  AND2 U39 (.A1(A[4]),.A2(B[5]),.Z(PP5[4]));
  AND2 U40 (.A1(A[5]),.A2(B[5]),.Z(PP5[5]));
  AND2 U41 (.A1(A[6]),.A2(B[5]),.Z(PP5[6]));
  AND2 u41 (.A1(A[7]),.A2(B[5]),.Z(PP5[7]));
  AND2 UU35 (.A1(A[8]),.A2(B[5]),.Z(PP5[8]));
  AND2 UU36 (.A1(A[9]),.A2(B[5]),.Z(PP5[9]));
  AND2 UU37 (.A1(A[10]),.A2(B[5]),.Z(PP5[10]));
  AND2 UU38 (.A1(A[11]),.A2(B[5]),.Z(PP5[11]));
  AND2 UU39 (.A1(A[12]),.A2(B[5]),.Z(PP5[12]));
  AND2 UU40 (.A1(A[13]),.A2(B[5]),.Z(PP5[13]));
  AND2 UU41 (.A1(A[14]),.A2(B[5]),.Z(PP5[14]));
  AND2 uU41 (.A1(A[15]),.A2(B[5]),.Z(PP5[15]));
////////////////// PP 6////////////////////////////
  AND2 U42 (.A1(A[0]),.A2(B[6]),.Z(PP6[0]));
  AND2 U43 (.A1(A[1]),.A2(B[6]),.Z(PP6[1]));
  AND2 U44 (.A1(A[2]),.A2(B[6]),.Z(PP6[2]));
  AND2 U45 (.A1(A[3]),.A2(B[6]),.Z(PP6[3]));
  AND2 U46 (.A1(A[4]),.A2(B[6]),.Z(PP6[4]));
  AND2 U47 (.A1(A[5]),.A2(B[6]),.Z(PP6[5]));
  AND2 U48 (.A1(A[6]),.A2(B[6]),.Z(PP6[6]));
  AND2 u48 (.A1(A[7]),.A2(B[6]),.Z(PP6[7]));
  AND2 UU42 (.A1(A[8]),.A2(B[6]),.Z(PP6[8]));
  AND2 UU43 (.A1(A[9]),.A2(B[6]),.Z(PP6[9]));
  AND2 UU44 (.A1(A[10]),.A2(B[6]),.Z(PP6[10]));
  AND2 UU45 (.A1(A[11]),.A2(B[6]),.Z(PP6[11]));
  AND2 UU46 (.A1(A[12]),.A2(B[6]),.Z(PP6[12]));
  AND2 UU47 (.A1(A[13]),.A2(B[6]),.Z(PP6[13]));
  AND2 UU48 (.A1(A[14]),.A2(B[6]),.Z(PP6[14]));
  AND2 uU48 (.A1(A[15]),.A2(B[6]),.Z(PP6[15]));
  ////////////////// PP 7////////////////////////////
  AND2 u49 (.A1(A[0]),.A2(B[7]),.Z(PP7[0]));
  AND2 u50 (.A1(A[1]),.A2(B[7]),.Z(PP7[1]));
  AND2 u51 (.A1(A[2]),.A2(B[7]),.Z(PP7[2]));
  AND2 u52 (.A1(A[3]),.A2(B[7]),.Z(PP7[3]));
  AND2 u53 (.A1(A[4]),.A2(B[7]),.Z(PP7[4]));
  AND2 u54 (.A1(A[5]),.A2(B[7]),.Z(PP7[5]));
  AND2 u55 (.A1(A[6]),.A2(B[7]),.Z(PP7[6]));
  AND2 u56 (.A1(A[7]),.A2(B[7]),.Z(PP7[7]));
  AND2 uU49 (.A1(A[8]),.A2(B[7]),.Z(PP7[8]));
  AND2 uU50 (.A1(A[9]),.A2(B[7]),.Z(PP7[9]));
  AND2 uU51 (.A1(A[10]),.A2(B[7]),.Z(PP7[10]));
  AND2 uU52 (.A1(A[11]),.A2(B[7]),.Z(PP7[11]));
  AND2 uU53 (.A1(A[12]),.A2(B[7]),.Z(PP7[12]));
  AND2 uU54 (.A1(A[13]),.A2(B[7]),.Z(PP7[13]));
  AND2 uU55 (.A1(A[14]),.A2(B[7]),.Z(PP7[14]));
  AND2 uU56 (.A1(A[15]),.A2(B[7]),.Z(PP7[15]));  
  ////////////////// PP 8 ////////////////////////////
  AND2 UX0 (.A1(A[0]),.A2(B[8]),.Z(PP8[0]));
  AND2 UX1 (.A1(A[1]),.A2(B[8]),.Z(PP8[1]));
  AND2 UX2 (.A1(A[2]),.A2(B[8]),.Z(PP8[2]));
  AND2 UX3 (.A1(A[3]),.A2(B[8]),.Z(PP8[3]));
  AND2 UX4 (.A1(A[4]),.A2(B[8]),.Z(PP8[4]));
  AND2 UX5 (.A1(A[5]),.A2(B[8]),.Z(PP8[5]));
  AND2 UX6 (.A1(A[6]),.A2(B[8]),.Z(PP8[6]));
  AND2 uX7 (.A1(A[7]),.A2(B[8]),.Z(PP8[7]));
  AND2 UXU0 (.A1(A[8]),.A2(B[8]),.Z(PP8[8]));
  AND2 UXU1 (.A1(A[9]),.A2(B[8]),.Z(PP8[9]));
  AND2 UXU2 (.A1(A[10]),.A2(B[8]),.Z(PP8[10]));
  AND2 UXU3 (.A1(A[11]),.A2(B[8]),.Z(PP8[11]));
  AND2 UXU4 (.A1(A[12]),.A2(B[8]),.Z(PP8[12]));
  AND2 UXU5 (.A1(A[13]),.A2(B[8]),.Z(PP8[13]));
  AND2 UXU6 (.A1(A[14]),.A2(B[8]),.Z(PP8[14]));
  AND2 uXU7 (.A1(A[15]),.A2(B[8]),.Z(PP8[15]));
////////////////// PP 9////////////////////////////
  AND2 UX7 (.A1(A[0]),.A2(B[9]),.Z(PP9[0]));
  AND2 UX8 (.A1(A[1]),.A2(B[9]),.Z(PP9[1]));
  AND2 UX9 (.A1(A[2]),.A2(B[9]),.Z(PP9[2]));
  AND2 UX10 (.A1(A[3]),.A2(B[9]),.Z(PP9[3]));
  AND2 UX11 (.A1(A[4]),.A2(B[9]),.Z(PP9[4]));
  AND2 UX12 (.A1(A[5]),.A2(B[9]),.Z(PP9[5]));
  AND2 UX13 (.A1(A[6]),.A2(B[9]),.Z(PP9[6]));
  AND2 uX14 (.A1(A[7]),.A2(B[9]),.Z(PP9[7]));
  AND2 UZU7 (.A1(A[8]),.A2(B[9]),.Z(PP9[8]));
  AND2 UXU8 (.A1(A[9]),.A2(B[9]),.Z(PP9[9]));
  AND2 UXU9 (.A1(A[10]),.A2(B[9]),.Z(PP9[10]));
  AND2 UXU10 (.A1(A[11]),.A2(B[9]),.Z(PP9[11]));
  AND2 UXU11 (.A1(A[12]),.A2(B[9]),.Z(PP9[12]));
  AND2 UXU12 (.A1(A[13]),.A2(B[9]),.Z(PP9[13]));
  AND2 UXU13 (.A1(A[14]),.A2(B[9]),.Z(PP9[14]));
  AND2 uXU14 (.A1(A[15]),.A2(B[9]),.Z(PP9[15]));
////////////////// PP 10////////////////////////////
  AND2 UX14 (.A1(A[0]),.A2(B[10]),.Z(PP10[0]));
  AND2 UX15 (.A1(A[1]),.A2(B[10]),.Z(PP10[1]));
  AND2 UX16 (.A1(A[2]),.A2(B[10]),.Z(PP10[2]));
  AND2 UX17 (.A1(A[3]),.A2(B[10]),.Z(PP10[3]));
  AND2 UX18 (.A1(A[4]),.A2(B[10]),.Z(PP10[4]));
  AND2 UX19 (.A1(A[5]),.A2(B[10]),.Z(PP10[5]));
  AND2 UX20 (.A1(A[6]),.A2(B[10]),.Z(PP10[6]));
  AND2 uX21 (.A1(A[7]),.A2(B[10]),.Z(PP10[7]));
  AND2 UZU14 (.A1(A[8]),.A2(B[10]),.Z(PP10[8]));
  AND2 UXU15 (.A1(A[9]),.A2(B[10]),.Z(PP10[9]));
  AND2 UXU16 (.A1(A[10]),.A2(B[10]),.Z(PP10[10]));
  AND2 UXU17 (.A1(A[11]),.A2(B[10]),.Z(PP10[11]));
  AND2 UXU18 (.A1(A[12]),.A2(B[10]),.Z(PP10[12]));
  AND2 UXU19 (.A1(A[13]),.A2(B[10]),.Z(PP10[13]));
  AND2 UXU20 (.A1(A[14]),.A2(B[10]),.Z(PP10[14]));
  AND2 UZu21 (.A1(A[15]),.A2(B[10]),.Z(PP10[15]));
////////////////// PP 11////////////////////////////
  AND2 UX21 (.A1(A[0]),.A2(B[11]),.Z(PP11[0]));
  AND2 UX22 (.A1(A[1]),.A2(B[11]),.Z(PP11[1]));
  AND2 UX23 (.A1(A[2]),.A2(B[11]),.Z(PP11[2]));
  AND2 UX24 (.A1(A[3]),.A2(B[11]),.Z(PP11[3]));
  AND2 UX25 (.A1(A[4]),.A2(B[11]),.Z(PP11[4]));
  AND2 UX26 (.A1(A[5]),.A2(B[11]),.Z(PP11[5]));
  AND2 UX27 (.A1(A[6]),.A2(B[11]),.Z(PP11[6]));
  AND2 uXU28 (.A1(A[7]),.A2(B[11]),.Z(PP11[7]));
  AND2 UXU21 (.A1(A[8]),.A2(B[11]),.Z(PP11[8]));
  AND2 UXU22 (.A1(A[9]),.A2(B[11]),.Z(PP11[9]));
  AND2 UXU23 (.A1(A[10]),.A2(B[11]),.Z(PP11[10]));
  AND2 UXU24 (.A1(A[11]),.A2(B[11]),.Z(PP11[11]));
  AND2 UXU25 (.A1(A[12]),.A2(B[11]),.Z(PP11[12]));
  AND2 UXU26 (.A1(A[13]),.A2(B[11]),.Z(PP11[13]));
  AND2 UXU27 (.A1(A[14]),.A2(B[11]),.Z(PP11[14]));
  AND2 UGU28 (.A1(A[15]),.A2(B[11]),.Z(PP11[15]));
////////X////////// PP 12////////////////////////////
  AND2 UX28 (.A1(A[0]),.A2(B[12]),.Z(PP12[0]));
  AND2 UX29 (.A1(A[1]),.A2(B[12]),.Z(PP12[1]));
  AND2 UX30 (.A1(A[2]),.A2(B[12]),.Z(PP12[2]));
  AND2 UX31 (.A1(A[3]),.A2(B[12]),.Z(PP12[3]));
  AND2 UX32 (.A1(A[4]),.A2(B[12]),.Z(PP12[4]));
  AND2 UX33 (.A1(A[5]),.A2(B[12]),.Z(PP12[5]));
  AND2 UX34 (.A1(A[6]),.A2(B[12]),.Z(PP12[6]));
  AND2 uX35 (.A1(A[7]),.A2(B[12]),.Z(PP12[7]));
  AND2 UZU28 (.A1(A[8]),.A2(B[12]),.Z(PP12[8]));
  AND2 UXU29 (.A1(A[9]),.A2(B[12]),.Z(PP12[9]));
  AND2 UXU30 (.A1(A[10]),.A2(B[12]),.Z(PP12[10]));
  AND2 UXU31 (.A1(A[11]),.A2(B[12]),.Z(PP12[11]));
  AND2 UXU32 (.A1(A[12]),.A2(B[12]),.Z(PP12[12]));
  AND2 UXU33 (.A1(A[13]),.A2(B[12]),.Z(PP12[13]));
  AND2 UXU34 (.A1(A[14]),.A2(B[12]),.Z(PP12[14]));
  AND2 uXR35 (.A1(A[15]),.A2(B[12]),.Z(PP12[15]));
////////X////////// PP 13////////////////////////////
  AND2 UX35 (.A1(A[0]),.A2(B[13]),.Z(PP13[0]));
  AND2 UX36 (.A1(A[1]),.A2(B[13]),.Z(PP13[1]));
  AND2 UX37 (.A1(A[2]),.A2(B[13]),.Z(PP13[2]));
  AND2 UX38 (.A1(A[3]),.A2(B[13]),.Z(PP13[3]));
  AND2 UX39 (.A1(A[4]),.A2(B[13]),.Z(PP13[4]));
  AND2 UX40 (.A1(A[5]),.A2(B[13]),.Z(PP13[5]));
  AND2 UX41 (.A1(A[6]),.A2(B[13]),.Z(PP13[6]));
  AND2 uX41 (.A1(A[7]),.A2(B[13]),.Z(PP13[7]));
  AND2 UXU35 (.A1(A[8]),.A2(B[13]),.Z(PP13[8]));
  AND2 UXU36 (.A1(A[9]),.A2(B[13]),.Z(PP13[9]));
  AND2 UXU37 (.A1(A[10]),.A2(B[13]),.Z(PP13[10]));
  AND2 UXU38 (.A1(A[11]),.A2(B[13]),.Z(PP13[11]));
  AND2 UXU39 (.A1(A[12]),.A2(B[13]),.Z(PP13[12]));
  AND2 UXU40 (.A1(A[13]),.A2(B[13]),.Z(PP13[13]));
  AND2 UZU41 (.A1(A[14]),.A2(B[13]),.Z(PP13[14]));
  AND2 uXU41 (.A1(A[15]),.A2(B[13]),.Z(PP13[15]));
////////X////////// PP 14////////////////////////////
  AND2 UX42 (.A1(A[0]),.A2(B[14]),.Z(PP14[0]));
  AND2 UX43 (.A1(A[1]),.A2(B[14]),.Z(PP14[1]));
  AND2 UX44 (.A1(A[2]),.A2(B[14]),.Z(PP14[2]));
  AND2 UX45 (.A1(A[3]),.A2(B[14]),.Z(PP14[3]));
  AND2 UX46 (.A1(A[4]),.A2(B[14]),.Z(PP14[4]));
  AND2 UX47 (.A1(A[5]),.A2(B[14]),.Z(PP14[5]));
  AND2 UX48 (.A1(A[6]),.A2(B[14]),.Z(PP14[6]));
  AND2 uX48 (.A1(A[7]),.A2(B[14]),.Z(PP14[7]));
  AND2 UXU42 (.A1(A[8]),.A2(B[14]),.Z(PP14[8]));
  AND2 UXU43 (.A1(A[9]),.A2(B[14]),.Z(PP14[9]));
  AND2 UXU44 (.A1(A[10]),.A2(B[14]),.Z(PP14[10]));
  AND2 UXU45 (.A1(A[11]),.A2(B[14]),.Z(PP14[11]));
  AND2 UXU46 (.A1(A[12]),.A2(B[14]),.Z(PP14[12]));
  AND2 UXU47 (.A1(A[13]),.A2(B[14]),.Z(PP14[13]));
  AND2 UXU48 (.A1(A[14]),.A2(B[14]),.Z(PP14[14]));
  AND2 XXU48 (.A1(A[15]),.A2(B[14]),.Z(PP14[15]));
  //////X//////////// PP 15////////////////////////////
  AND2 uX49 (.A1(A[0]),.A2(B[15]),.Z(PP15[0]));
  AND2 uX50 (.A1(A[1]),.A2(B[15]),.Z(PP15[1]));
  AND2 uX51 (.A1(A[2]),.A2(B[15]),.Z(PP15[2]));
  AND2 uX52 (.A1(A[3]),.A2(B[15]),.Z(PP15[3]));
  AND2 uX53 (.A1(A[4]),.A2(B[15]),.Z(PP15[4]));
  AND2 uX54 (.A1(A[5]),.A2(B[15]),.Z(PP15[5]));
  AND2 uX55 (.A1(A[6]),.A2(B[15]),.Z(PP15[6]));
  AND2 uX56 (.A1(A[7]),.A2(B[15]),.Z(PP15[7]));
  AND2 uXU49 (.A1(A[8]),.A2(B[15]),.Z(PP15[8]));
  AND2 uXU50 (.A1(A[9]),.A2(B[15]),.Z(PP15[9]));
  AND2 uXU51 (.A1(A[10]),.A2(B[15]),.Z(PP15[10]));
  AND2 uXU52 (.A1(A[11]),.A2(B[15]),.Z(PP15[11]));
  AND2 uXU53 (.A1(A[12]),.A2(B[15]),.Z(PP15[12]));
  AND2 uXU54 (.A1(A[13]),.A2(B[15]),.Z(PP15[13]));
  AND2 uXU55 (.A1(A[14]),.A2(B[15]),.Z(PP15[14]));
  AND2 uXU56 (.A1(A[15]),.A2(B[15]),.Z(PP15[15])); 
  
  endmodule